//pwm module, outputs a pulse width according to the value written
//max width 255 cycles

module pwm(input clk, input en, input [7:0] value_input, output out);

   
endmodule
